`include "..\maraudersv\marauder.sv"

module regstb(
    
);

endmodule